`define SSC_IFID 4
`define SSC_IX   4
`define SSC_IL   1
`define SSC_IS   1

`define MEM_RPORTS (`SSC_IFID + `SSC_IL)
