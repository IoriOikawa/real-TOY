`define SSC_IF (`SSC_EX)
`define SSC_EX 5
`define SSC_MEM 1 // fixed

`define MEM_RPORTS (`SSC_IF)

`define I2C_DIV 192 // 12MHz -> 62.5kHz
