`include "global.svh"

interface core_arf_r;
   logic [3:0] addr;
   logic [15:0] data;
endinterface
