`define SSC_IF (`SSC_EX + `SSC_MEM)
`define SSC_EX 5
`define SSC_MEM 1

`define MEM_RPORTS (`SSC_IF)
